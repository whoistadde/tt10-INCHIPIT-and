//  Module: and_module
//

module and_module
    (
        input logic a,
        input logic b,
        output logic y
    );

    assign y = a & b;
endmodule: and_module
